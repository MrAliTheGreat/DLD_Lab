library verilog;
use verilog.vl_types.all;
entity AlternativeTB is
end AlternativeTB;
